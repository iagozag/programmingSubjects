`ifndef DEFINITIONS_SV
`define DEFINITIONS_SV

// Definições globais da mensagem a ser encriptada
`define MSG_SIZE 128
`define MSG 128'b0011011101010110100101111100110001101100100100011101000101101101111011011101101001001100100011011001101010101110000101011001110

`endif

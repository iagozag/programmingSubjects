`include "definitions.sv"
`include "shifter.sv"
`include "cypher.sv"
